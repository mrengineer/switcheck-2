`timescale 1 ns / 1 ps

module ADC #
(
  parameter integer ADC_DATA_WIDTH = 14
)
(
  // System signals
  input  wire        aclk,
  input  wire        aresetn,      // Active-low reset

  // ADC signals
  output wire        adc_csn,
  input  wire [15:0] adc_dat_a,
  input  wire [15:0] adc_dat_b,

  output wire [15:0] cur_adc,
  output wire [63:0] cur_sample,
  
  input wire  [7:0] limiter,           // Сколько писать отсчетов в серии максимум (число 2^limiter) 
  


  // Trigger level setting
  input  wire [15:0] trigger_level,

  // Reset control signals
  input  wire        reset_trigger,     // Сброс триггера при 1 извне
  input  wire        reset_max_sum,     // Сброс максимума суммы при 1

  // AXI-Stream master (32-bit words)
  output reg         m_axis_tvalid,
  output wire [31:0] m_axis_tdata,
  
  // Output for max_sum_abs
  output reg  signed [15:0] max_sum_out,
  output reg  [63:0]        last_detrigged,     // последний раз пересекли триггер вниз
  output reg  [63:0]        first_trigged,      // первый раз сработал триггер
  output reg  [63:0]        cur_limiter,        // Ограничивает запись числом записей на одну серию
  output reg  [31:0]        samples_sent,       // Число отсчётов, сохранённых в шину
  output reg                trigger_activated,  // Флаг активации триггера
  output reg  [15:0]        triggers_count      // сколько раз сработал триггер
);

  // =========================
  // Параметры и внутренности
  // =========================

  localparam PADDING_WIDTH = 16 - ADC_DATA_WIDTH;
  localparam MID_SCALE     = 1 << (ADC_DATA_WIDTH-1); // для 14 бит: 0x2000
 

  // Сырые/обработанные данные
  reg  signed [ADC_DATA_WIDTH-1:0] int_dat_a_reg; // signed
  reg  signed [ADC_DATA_WIDTH-1:0] int_dat_b_reg; // signed
  reg         [ADC_DATA_WIDTH-1:0] abs_a;
  reg         [ADC_DATA_WIDTH-1:0] abs_b;
  reg         [ADC_DATA_WIDTH:0]   sum_abs;       // +1 бит на сумму
  reg         [15:0]               max_sum_abs;

  reg  [63:0] sample_counter;

  // =========================
  // Формирование AXI-выхода
  // =========================

  reg [31:0] axis_data_reg;   // Регистр данных на выход
  assign m_axis_tdata = axis_data_reg;

  // Флаги событий для посылки служебных пакетов
  reg prev_trigger_activated;
  reg need_send_cnt_low;
  reg need_send_cnt_high;
  reg need_send_end;


  wire [63:0] limiter_val;             // чтобы ограничить limiter, 
  // ограничиваем максимум 63, иначе будет переполнение при (1 << limiter)
  assign limiter_val = (limiter > 8'd63) ? 64'hFFFF_FFFF_FFFF_FFFF : (64'd1 << limiter);


  // =========================
  // Подготовка 15-бит unsigned A/B
  // =========================
  // Сместим signed к unsigned и ограничим в 0..32767 (15 бит).
  // Для корректности на любой ADC_DATA_WIDTH<=15.
  wire signed [15:0] a_ext = {{(16-ADC_DATA_WIDTH){int_dat_a_reg[ADC_DATA_WIDTH-1]}}, int_dat_a_reg};
  wire signed [15:0] b_ext = {{(16-ADC_DATA_WIDTH){int_dat_b_reg[ADC_DATA_WIDTH-1]}}, int_dat_b_reg};

  // Берём 15 младших бит, со знаком
  wire [14:0] a_u15 = a_ext[14:0];
  wire [14:0] b_u15 = b_ext[14:0];


  // =========================
  // Основной процесс
  // =========================

  always @(posedge aclk or negedge aresetn) begin
    if (!aresetn) begin
      int_dat_a_reg         <= 0;
      int_dat_b_reg         <= 0;
      abs_a                 <= 0;
      abs_b                 <= 0;
      sum_abs               <= 0;
      m_axis_tvalid         <= 1'b0;
      axis_data_reg         <= 32'd0;

      trigger_activated     <= 1'b0;
      prev_trigger_activated<= 1'b0;
      triggers_count        <= 0;
      max_sum_abs           <= 0;
      sample_counter        <= 64'd0;
      samples_sent          <= 0;
      max_sum_out           <= 0;
      last_detrigged        <= 0;
      first_trigged         <= 0;
      cur_limiter           <= 0;

      need_send_cnt_low     <= 1'b0;
      need_send_cnt_high    <= 1'b0;
      need_send_end         <= 1'b0;

    end else begin

      // -------------------------
      // Сброс части триггера
      // -------------------------
      if (reset_trigger) begin
        last_detrigged        <= 0;
        first_trigged         <= 0;
        triggers_count        <= 0;
        trigger_activated     <= 1'b1;      //  временно 1!
        cur_limiter           <= 0;
        need_send_end         <= 1'b0;
        need_send_cnt_low     <= 1'b0;
        need_send_cnt_high    <= 1'b0;
        
        
        sample_counter <= 64'd0;                //временно!
      end


      last_detrigged <= limiter;

      // -------------------------
      // Счётчик семплов
      // -------------------------
      sample_counter <= sample_counter + 1;

      // -------------------------
      // Захват и нормализация ADC
      // (адаптировано из исходника)
      // -------------------------
      int_dat_a_reg <= {{(PADDING_WIDTH+1){adc_dat_a[ADC_DATA_WIDTH-1]}}, ~adc_dat_a[ADC_DATA_WIDTH-2:0]} + MID_SCALE;
      int_dat_b_reg <= {{(PADDING_WIDTH+1){adc_dat_b[ADC_DATA_WIDTH-1]}}, ~adc_dat_b[ADC_DATA_WIDTH-2:0]} + MID_SCALE;

      abs_a <= int_dat_a_reg[ADC_DATA_WIDTH-1] ? (~int_dat_a_reg + 1) : int_dat_a_reg;
      abs_b <= int_dat_b_reg[ADC_DATA_WIDTH-1] ? (~int_dat_b_reg + 1) : int_dat_b_reg;

      sum_abs <= abs_a + abs_b;

        // Трекинг максимума
        if (sum_abs > max_sum_abs && !reset_max_sum)
          max_sum_abs <= sum_abs;
        else if (reset_max_sum)
          max_sum_abs <= 0;

        // -------------------------
        // Логика триггера
        // -------------------------
        // Включение
        /*if (sum_abs > trigger_level && !reset_trigger && trigger_activated == 1'b0) begin
          cur_limiter           <= 0;
          first_trigged         <= sample_counter;
          trigger_activated     <= 1'b1;
          triggers_count        <= triggers_count + 1;

          // При фронте триггера нужно отправить счётчик (2 слова)
          need_send_cnt_low     <= 1'b1;
          need_send_cnt_high    <= 1'b1;
        end*/

        // Выключение (по уровню)
        /*
        if (sum_abs < trigger_level && !reset_trigger && trigger_activated == 1'b1) begin
          last_detrigged        <= sample_counter;
          trigger_activated     <= 1'b0;
          need_send_end         <= 1'b1;   // по спаду - отправить окончание
        end
        */



        // Ограничение длины серии
        //if (cur_limiter > limiter*10 && trigger_activated == 1'b1) begin
        /*if (cur_limiter >= limiter_val && trigger_activated == 1'b1) begin
          trigger_activated     <= 1'b0;   // отрубить
          need_send_end         <= 1'b1;   // и отправить окончание
        end*/


        // Вывод статистики
        max_sum_out <= max_sum_abs;

      // -------------------------
      // Формирование AXI-Stream
      // Очерёдность: cnt_low -> cnt_high -> data(если активен) -> end
      // За такт уходит максимум 1 слово.
      // -------------------------
      m_axis_tvalid <= 1'b0; // по умолчанию



      //if (sample_counter < 64'd150) begin   // Временно

      // Фронт/спад триггера детектируем
      prev_trigger_activated <= trigger_activated;

      // 1) Если нужно отправить счетчик (после фронта)
      /*if (need_send_cnt_low) begin
        axis_data_reg     <= {2'b00, sample_counter[29:0]};
        m_axis_tvalid     <= 1'b1;
        need_send_cnt_low <= 1'b0;
      end else if (need_send_cnt_high) begin
        axis_data_reg      <= {2'b01, sample_counter[59:30]};
        m_axis_tvalid      <= 1'b1;
        need_send_cnt_high <= 1'b0;

      // 2) Пока активен триггер - шлём данные АЦП
      end else */
      
      if (trigger_activated) begin       
        cur_limiter           <= cur_limiter + 1;
        samples_sent          <= samples_sent + 1;
                  
        axis_data_reg  <= {2'b10, 15'd123, 15'd555};
        m_axis_tvalid  <= 1'b1;
        
        if (samples_sent > 32'd32) begin 
            trigger_activated  <= 1'b0;
        end               
      end

      /*
      // 3) Если нужно отправить окончание
      end else if (need_send_end) begin
        axis_data_reg  <= {2'b11, 30'd0};
        m_axis_tvalid  <= 1'b1;
        need_send_end  <= 1'b0;
      end
      */
      
      
      //end
      
    end
  end




  // =========================
  // Прочие связи
  // =========================

  assign adc_csn     = 1'b1;
  assign cur_adc     = sum_abs;
  assign cur_sample  = sample_counter;

endmodule

